`timescale 1ns / 1ps

module invroundlast(
    input [3:0]rc,
    input [127:0]data,
    input [127:0]keylastin,
    output [127:0]fout
);

wire [127:0] sb,sr,mcl,keyout;

invKeyGeneration t0(rc,keylastin,keyout);
invshiftrow t2(data,sr);
invsubbytes t1(sr,sb);
assign fout= keyout^sb;

endmodule
