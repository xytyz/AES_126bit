`timescale 1ns / 1ps

module invsbox(
input  [7:0] a,
output reg [7:0] c);
    
    
   always @(a)
    case (a)
        8'h00: c = 8'h52;
        8'h01: c = 8'h09;
        8'h02: c = 8'h6A;
        8'h03: c = 8'hD5;
        8'h04: c = 8'h30;
        8'h05: c = 8'h36;
        8'h06: c = 8'hA5;
        8'h07: c = 8'h38;
        8'h08: c = 8'hBF;
        8'h09: c = 8'h40;
        8'h0A: c = 8'hA3;
        8'h0B: c = 8'h9E;
        8'h0C: c = 8'h81;
        8'h0D: c = 8'hF3;
        8'h0E: c = 8'hD7;
        8'h0F: c = 8'hFB;
        8'h10: c = 8'h7C;
        8'h11: c = 8'hE3;
        8'h12: c = 8'h39;
        8'h13: c = 8'h82;
        8'h14: c = 8'h9B;
        8'h15: c = 8'h2F;
        8'h16: c = 8'hFF;
        8'h17: c = 8'h87;
        8'h18: c = 8'h34;
        8'h19: c = 8'h8E;
        8'h1A: c = 8'h43;
        8'h1B: c = 8'h44;
        8'h1C: c = 8'hC4;
        8'h1D: c = 8'hDE;
        8'h1E: c = 8'hE9;
        8'h1F: c = 8'hCB;
        8'h20: c = 8'h54;
        8'h21: c = 8'h7B;
        8'h22: c = 8'h94;
        8'h23: c = 8'h32;
        8'h24: c = 8'hA6;
        8'h25: c = 8'hC2;
        8'h26: c = 8'h23;
        8'h27: c = 8'h3D;
        8'h28: c = 8'hEE;
        8'h29: c = 8'h4C;
        8'h2A: c = 8'h95;
        8'h2B: c = 8'h0B;
        8'h2C: c = 8'h42;
        8'h2D: c = 8'hFA;
        8'h2E: c = 8'hC3;
        8'h2F: c = 8'h4E;
        8'h30: c = 8'h08;
        8'h31: c = 8'h2E;
        8'h32: c = 8'hA1;
        8'h33: c = 8'h66;
        8'h34: c = 8'h28;
        8'h35: c = 8'hD9;
        8'h36: c = 8'h24;
        8'h37: c = 8'hB2;
        8'h38: c = 8'h76;
        8'h39: c = 8'h5B;
        8'h3A: c = 8'hA2;
        8'h3B: c = 8'h49;
        8'h3C: c = 8'h6D;
        8'h3D: c = 8'h8B;
        8'h3E: c = 8'hD1;
        8'h3F: c = 8'h25;
        8'h40: c = 8'h72;
        8'h41: c = 8'hF8;
        8'h42: c = 8'hF6;
        8'h43: c = 8'h64;
        8'h44: c = 8'h86;
        8'h45: c = 8'h68;
        8'h46: c = 8'h98;
        8'h47: c = 8'h16;
        8'h48: c = 8'hD4;
        8'h49: c = 8'hA4;
        8'h4A: c = 8'h5C;
        8'h4B: c = 8'hCC;
        8'h4C: c = 8'h5D;
        8'h4D: c = 8'h65;
        8'h4E: c = 8'hB6;
        8'h4F: c = 8'h92;
        8'h50: c = 8'h6C;
        8'h51: c = 8'h70;
        8'h52: c = 8'h48;
        8'h53: c = 8'h50;
        8'h54: c = 8'hFD;
        8'h55: c = 8'hED;
        8'h56: c = 8'hB9;
        8'h57: c = 8'hDA;
        8'h58: c = 8'h5E;
        8'h59: c = 8'h15;
        8'h5A: c = 8'h46;
        8'h5B: c = 8'h57;
        8'h5C: c = 8'hA7;
        8'h5D: c = 8'h8D;
        8'h5E: c = 8'h9D;
        8'h5F: c = 8'h84;
        8'h60: c = 8'h90;
        8'h61: c = 8'hD8;
        8'h62: c = 8'hAB;
        8'h63: c = 8'h00;
        8'h64: c = 8'h8C;
        8'h65: c = 8'hBC;
        8'h66: c = 8'hD3;
        8'h67: c = 8'h0A;
        8'h68: c = 8'hF7;
        8'h69: c = 8'hE4;
        8'h6A: c = 8'h58;
        8'h6B: c = 8'h05;
        8'h6C: c = 8'hB8;
        8'h6D: c = 8'hB3;
        8'h6E: c = 8'h45;
        8'h6F: c = 8'h06;
        8'h70: c = 8'hD0;
        8'h71: c = 8'h2C;
        8'h72: c = 8'h1E;
        8'h73: c = 8'h8F;
        8'h74: c = 8'hCA;
        8'h75: c = 8'h3F;
        8'h76: c = 8'h0F;
        8'h77: c = 8'h02;
        8'h78: c = 8'hC1;
        8'h79: c = 8'hAF;
        8'h7A: c = 8'hBD;
        8'h7B: c = 8'h03;
        8'h7C: c = 8'h01;
        8'h7D: c = 8'h13;
        8'h7E: c = 8'h8A;
        8'h7F: c = 8'h6B;
        8'h80: c = 8'h3A;
        8'h81: c = 8'h91;
        8'h82: c = 8'h11;
        8'h83: c = 8'h41;
        8'h84: c = 8'h4F;
        8'h85: c = 8'h67;
        8'h86: c = 8'hDC;
        8'h87: c = 8'hEA;
        8'h88: c = 8'h97;
        8'h89: c = 8'hF2;
        8'h8A: c = 8'hCF;
        8'h8B: c = 8'hCE;
        8'h8C: c = 8'hF0;
        8'h8D: c = 8'hB4;
        8'h8E: c = 8'hE6;
        8'h8F: c = 8'h73;
        8'h90: c = 8'h96;
        8'h91: c = 8'hAC;
        8'h92: c = 8'h74;
        8'h93: c = 8'h22;
        8'h94: c = 8'hE7;
        8'h95: c = 8'hAD;
        8'h96: c = 8'h35;
        8'h97: c = 8'h85;
        8'h98: c = 8'hE2;
        8'h99: c = 8'hF9;
        8'h9A: c = 8'h37;
        8'h9B: c = 8'hE8;
        8'h9C: c = 8'h1C;
        8'h9D: c = 8'h75;
        8'h9E: c = 8'hDF;
        8'h9F: c = 8'h6E;
        8'hA0: c = 8'h47;
        8'hA1: c = 8'hF1;
        8'hA2: c = 8'h1A;
        8'hA3: c = 8'h71;
        8'hA4: c = 8'h1D;
        8'hA5: c = 8'h29;
        8'hA6: c = 8'hC5;
        8'hA7: c = 8'h89;
        8'hA8: c = 8'h6F;
        8'hA9: c = 8'hB7;
        8'hAA: c = 8'h62;
        8'hAB: c = 8'h0E;
        8'hAC: c = 8'hAA;
        8'hAD: c = 8'h18;
        8'hAE: c = 8'hBE;
        8'hAF: c = 8'h1B;
        8'hB0: c = 8'hFC;
        8'hB1: c = 8'h56;
        8'hB2: c = 8'h3E;
        8'hB3: c = 8'h4B;
        8'hB4: c = 8'hC6;
        8'hB5: c = 8'hD2;
        8'hB6: c = 8'h79;
        8'hB7: c = 8'h20;
        8'hB8: c = 8'h9A;
        8'hB9: c = 8'hDB;
        8'hBA: c = 8'hC0;
        8'hBB: c = 8'hFE;
        8'hBC: c = 8'h78;
        8'hBD: c = 8'hCD;
        8'hBE: c = 8'h5A;
        8'hBF: c = 8'hF4;
        8'hC0: c = 8'h1F;
        8'hC1: c = 8'hDD;
        8'hC2: c = 8'hA8;
        8'hC3: c = 8'h33;
        8'hC4: c = 8'h88;
        8'hC5: c = 8'h07;
        8'hC6: c = 8'hC7;
        8'hC7: c = 8'h31;
        8'hC8: c = 8'hB1;
        8'hC9: c = 8'h12;
        8'hCA: c = 8'h10;
        8'hCB: c = 8'h59;
        8'hCC: c = 8'h27;
        8'hCD: c = 8'h80;
        8'hCE: c = 8'hEC;
        8'hCF: c = 8'h5F;
        8'hD0: c = 8'h60;
        8'hD1: c = 8'h51;
        8'hD2: c = 8'h7F;
        8'hD3: c = 8'hA9;
        8'hD4: c = 8'h19;
        8'hD5: c = 8'hB5;
        8'hD6: c = 8'h4A;
        8'hD7: c = 8'h0D;
        8'hD8: c = 8'h2D;
        8'hD9: c = 8'hE5;
        8'hDA: c = 8'h7A;
        8'hDB: c = 8'h9F;
        8'hDC: c = 8'h93;
        8'hDD: c = 8'hC9;
        8'hDE: c = 8'h9C;
        8'hDF: c = 8'hEF;
        8'hE0: c = 8'hA0;
        8'hE1: c = 8'hE0;
        8'hE2: c = 8'h3B;
        8'hE3: c = 8'h4D;
        8'hE4: c = 8'hAE;
        8'hE5: c = 8'h2A;
        8'hE6: c = 8'hF5;
        8'hE7: c = 8'hB0;
        8'hE8: c = 8'hC8;
        8'hE9: c = 8'hEB;
        8'hEA: c = 8'hBB;
        8'hEB: c = 8'h3C;
        8'hEC: c = 8'h83;
        8'hED: c = 8'h53;
        8'hEE: c = 8'h99;
        8'hEF: c = 8'h61;
        8'hF0: c = 8'h17;
        8'hF1: c = 8'h2B;
        8'hF2: c = 8'h04;
        8'hF3: c = 8'h7E;
        8'hF4: c = 8'hBA;
        8'hF5: c = 8'h77;
        8'hF6: c = 8'hD6;
        8'hF7: c = 8'h26;
        8'hF8: c = 8'hE1;
        8'hF9: c = 8'h69;
        8'hFA: c = 8'h14;
        8'hFB: c = 8'h63;
        8'hFC: c = 8'h55;
        8'hFD: c = 8'h21;
        8'hFE: c = 8'h0C;
        8'hFF: c = 8'h7D;
	endcase

endmodule
